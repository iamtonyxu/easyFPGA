module adder(  
    input   [3:0] a,  // First 4-bit input  
    input   [3:0] b,  // Second 4-bit input  
    input         cin, // Carry-in  
    output  [3:0] s,  // 4-bit sum  
    output        cout  // Carry-out  
);  


// Calculate each bit of the sum and carry  
// Using bitwise XOR for sum and AND for carry  
assign s[0] = a[0] ^ b[0] ^ cin;  
assign s[1] = a[1] ^ b[1] ^ (a[0] & b[0]);  
assign s[2] = a[2] ^ b[2] ^ (a[1] & b[1]);  
assign s[3] = a[3] ^ b[3] ^ (a[2] & b[2]);  

// The final carry-out is generated by the most significant bit addition  
assign cout = a[3] & b[3] | (a[2] & b[2]) | (a[1] & b[1]) | (a[0] & b[0]);  


//assign {cout, s} = a + b + cin;

endmodule